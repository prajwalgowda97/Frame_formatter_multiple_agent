package frame_formatter_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  // Sequence
  `include "./../uvme/sequences/frame_formatter_fifo_seq_item.sv"
  `include "./../uvme/sequences/frame_formatter_packet_seq_item.sv"
  `include "./../uvme/sequences/frame_formatter_header_seq_item.sv"
  `include "./../uvme/sequences/frame_formatter_fifo_sequence.sv"
  `include "./../uvme/sequences/frame_formatter_packet_sequence.sv"
  `include "./../uvme/sequences/frame_formatter_header_sequence.sv"
 




  // fifo agent 
  
  
    `include "./../uvme/fifoagent/frame_formatter_fifo_seqr.sv"
  `include "./../uvme/fifoagent/frame_formatter_fifo_driver.sv"
  `include "./../uvme/fifoagent/frame_formatter_fifo_monitor.sv"
  `include "./../uvme/fifoagent/frame_formatter_fifo_agent.sv"


  // packet agent
  `include "./../uvme/packetagent/frame_formatter_packet_seqr.sv"
   `include "./../uvme/packetagent/frame_formatter_packet_driver.sv"
  `include "./../uvme/packetagent/frame_formatter_packet_monitor.sv"
  `include "./../uvme/packetagent/frame_formatter_packet_agent.sv"


  // header agent
    `include "./../uvme/headeragent/frame_formatter_header_seqr.sv"
   `include "./../uvme/headeragent/frame_formatter_header_driver.sv"
  `include "./../uvme/headeragent/frame_formatter_header_monitor.sv"
  `include "./../uvme/headeragent/frame_formatter_header_agent.sv"


  // Enviornment
  `include "./../uvme/env/frame_formatter_coverage_model.sv"
  `include "./../uvme/env/frame_formatter_scoreboard.sv"
  `include "./../uvme/env/frame_formatter_env.sv"



  // test
  // Test
// `include "./../uvme/test/frame_formatter_base_test.sv"
 `include "./../uvme/test/frame_formatter_initial_reset_test.sv"
`include "./../uvme/test/frame_formatter_soft_reset_test.sv"
 `include "./../uvme/test/frame_formatter_reset_scenarios_test.sv"
`include "./../uvme/test/frame_formatter_ibypass_enable_test.sv"
 `include "./../uvme/test/frame_formatter_ibypass_disable_test.sv"
`include "./../uvme/test/frame_formatter_sync_fifo_full_test.sv"
`include "./../uvme/test/frame_formatter_async_fifo_empty_test.sv"
`include "./../uvme/test/frame_formatter_vlan_tag_disable_test.sv"
`include "./../uvme/test/frame_formatter_multiple_write_multiple_read_test.sv"
`include "./../uvme/test/frame_formatter_multiple_write_one_read_test.sv"
`include "./../uvme/test/frame_formatter_zero_write_multiple_read_test.sv"
`include "./../uvme/test/frame_formatter_random_write_read_test.sv"
`include "./../uvme/test/frame_formatter_ibypass_vlan_random_test.sv"












 endpackage
