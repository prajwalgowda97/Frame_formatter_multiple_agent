interface frame_formatter_clk_interface();

	logic Frame_Formatter_TOP_clk;
	logic async_fifo_rd_clk;

endinterface
